`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/07/2022 09:27:39 PM
// Design Name: 
// Module Name: Sim_Comp_Signed_4Bit
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Sim_Comp_Signed_4Bit(
      );
      
      // INPUTS
      reg A3;
      reg A2;
      reg A1;
      reg A0;
      reg B3;
      reg B2;
      reg B1;
      reg B0;
      
      // OUTPUTS
      wire A_GREATER_B;
      wire A_LESS_B;
      wire A_EQUAL_B;
     
      
      Comparator_Signed_4Bit UUT (
      .A3(A3),
      .A2(A2),
      .A1(A1),
      .A0(A0),
      
      .B3(B3),
      .B2(B2),
      .B1(B1),
      .B0(B0),
      
      .A_GREATER_B(A_GREATER_B),
      .A_LESS_B(A_LESS_B),
      .A_EQUAL_B(A_EQUAL_B)
      );
      
      // INITIALIZE INPUTS
      initial begin
          // --------------------------------------
          // TEST #1 
          // A = 0 // B = -8
          // --------------------------------------
          A3 = 0;
          A2 = 0;
          A1 = 0;
          A0 = 0;
          
          B3 = 1;
          B2 = 0;
          B1 = 0;
          B0 = 0;
          #10;
          
          // --------------------------------------
          // TEST #2
          // A = -8 // B = -1
          // --------------------------------------
          A3 = 1;
          A2 = 0;
          A1 = 0;
          A0 = 0;
            
          B3 = 1;
          B2 = 1;
          B1 = 1;
          B0 = 1;
          #10;
          
          // --------------------------------------
          // TEST #3
          // A = +7 // B = +3
          // --------------------------------------
          A3 = 0;
          A2 = 1;
          A1 = 1;
          A0 = 1;
            
          B3 = 0;
          B2 = 0;
          B1 = 1;
          B0 = 1;
          #10;
          
          // --------------------------------------
          // TEST #4
          // A = -7 // B = +1
          // --------------------------------------
          A3 = 1;
          A2 = 0;
          A1 = 0;
          A0 = 1;
            
          B3 = 0;
          B2 = 0;
          B1 = 0;
          B0 = 1;
          #10;
          
          // --------------------------------------
          // TEST #5
          // A = +4 // B = -4
          // --------------------------------------
          A3 = 0;
          A2 = 1;
          A1 = 0;
          A0 = 0;
            
          B3 = 1;
          B2 = 1;
          B1 = 0;
          B0 = 0;
          #10;
          
          // --------------------------------------
          // TEST #6
          // A = -2 // B = -2
          // --------------------------------------
          A3 = 1;
          A2 = 1;
          A1 = 1;
          A0 = 0;
            
          B3 = 1;
          B2 = 1;
          B1 = 1;
          B0 = 0;
          #10;
          
          // --------------------------------------
          // TEST #7
          // A = 5 // B = 2
          // --------------------------------------
          A3 = 0;
          A2 = 1;
          A1 = 0;
          A0 = 0;
            
          B3 = 0;
          B2 = 0;
          B1 = 1;
          B0 = 0;
          #10;
          
          // --------------------------------------
          // TEST #8
          // A = -1 // B = -1
          // --------------------------------------
          A3 = 1;
          A2 = 1;
          A1 = 1;
          A0 = 1;
            
          B3 = 1;
          B2 = 1;
          B1 = 1;
          B0 = 1;
          #10;
         
      end 
endmodule
